`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:13:28 12/09/2013 
// Design Name: 
// Module Name:    iqdemap_bpsk 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module iqmap_qpsk(
    input CLK,
    input RST,
    input ce,
    input valid_i,
    input [127:0] input,
    input reader_en,
    output [10:0] xr,
    output [10:0] xi,
    output valid_o,
    output valid_raw,
    output [3:0] raw
    );


endmodule
