`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:18:14 12/09/2013 
// Design Name: 
// Module Name:    iqdemap_bpsk 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module iqdemap_bpsk(
                    input               CLK,
                    input               RST,
                    input               ce,
                    input               valid_i,
                    input signed [10:0] ar,
                    input signed [10:0] ai,
                    output reg          valid_o,
                    output reg [127:0]  writer_data,
                    output              valid_raw,
                    output reg [3:0]    raw
                    );

   reg [8:0]                            cnt;
   reg                                  write_data_output_flg;

   assign valid_raw = valid_o;
   
   
   always@(posedge CLK)
     begin
        if(!RST)
          begin
             cnt <= 0;
             
             valid_o <= 0;
             raw <= 0;
          end
        else
          begin
             if(write_data_output_flg)  
               begin
                  cnt <= 0;
                  write_data_output_flg <= 0;
                  valid_o <= 0;              
               end
             else
               begin
                  if(valid_i)
                    begin
                       raw <= ar;
                       writer_data[cnt] <= ((1 - ar) >> 1);
                       cnt <= cnt + 1;
                       if(cnt >= 128)
                         begin
                            write_data_output_flg <= 1;
                            valid_o <= 1;
                         end
                    end
                  else
                    begin
                       cnt <= 0;
                    end 
               end 
          end
        
     end
   

   
endmodule
